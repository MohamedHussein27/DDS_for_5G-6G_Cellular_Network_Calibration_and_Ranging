// this package has the shared signals among packages
package alu_shared_pkg;
    // counters
    int error_count_out = 0; 
    int correct_count_out = 0;
    int error_count_c = 0;
    int correct_count_c = 0;
endpackage