package shared_pkg;
    typedef enum  {
            IDLE    ,
            S1      ,
            S10     ,
            S101    
        } state_e; 
    state_e cs, ns;
endpackage

