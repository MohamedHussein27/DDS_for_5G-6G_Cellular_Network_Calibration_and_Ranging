package alu_pack;

typedef enum {ADD_op=0, XOR_op=1, AND_op=2, OR_op=3} operation_t;
    
endpackage