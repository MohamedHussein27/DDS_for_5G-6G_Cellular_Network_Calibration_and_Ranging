package alu_pkg;

  typedef enum bit [1:0] {
    ADD_op=0,
     XOR_op=1,
      AND_op=2,
       OR_op=3
  } opcode_t;


    
endpackage