// this package has the shared signals among packages
package shared_pkg;
    int test_finished; // when high, stop the simulation
    // counters
    int error_count_out = 0; 
    int correct_count_out = 0;
    int error_count_c = 0;
    int correct_count_c = 0;
endpackage