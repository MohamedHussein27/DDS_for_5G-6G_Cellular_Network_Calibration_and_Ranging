package alu_scoreboard_pkg;
    import alu_seq_item_pkg::*;
    import shared_pkg::*;
    class alu_scoreboard;
        
        // reference signals
        logic [3:0] out_ref;
        logic c_ref;

        // compare function
        function void check_data (alu_seq_item tr);
            reference_model(tr);
            // compare
            if (tr.out !== out_ref) begin
                error_count_out++;
                $display("error in data out, ref_out is: %0d     while dut out is: %0d", out_ref, tr.out);
            end
            else
                correct_count_out++;
            if(tr.c !== c_ref) begin
                error_count_c++;
                $display("error in carry, ref_c is: %0d    while dut c is: %0d", c_ref, tr.c);
            end
            else
                correct_count_c++;
        endfunction
        // reference function
        function void reference_model (alu_seq_item tr_ref);
            case (tr_ref.op)
                2'b00: begin // addition
                    {c_ref, out_ref} = tr_ref.a + tr_ref.b;
                end
                2'b01: begin // XOR
                    c_ref = 0;
                    out_ref = tr_ref.a ^ tr_ref.b;
                end
                2'b10: begin // AND
                    c_ref = 0;
                    out_ref = tr_ref.a &  tr_ref.b;
                end
                2'b11: begin // OR
                    c_ref = 0;
                    out_ref = tr_ref.a | tr_ref.b;
                end
                default: begin
                    c_ref = 0;
                    out_ref = 4'b0000;
                end
            endcase
        endfunction
    endclass
endpackage